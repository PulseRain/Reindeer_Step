/*
###############################################################################
# Copyright (c) 2019, PulseRain Technology LLC 
#
# This program is distributed under a dual license: an open source license, 
# and a commercial license. 
# 
# The open source license under which this program is distributed is the 
# GNU Public License version 3 (GPLv3).
#
# And for those who want to use this program in ways that are incompatible
# with the GPLv3, PulseRain Technology LLC offers commercial license instead.
# Please contact PulseRain Technology LLC (www.pulserain.com) for more detail.
#
###############################################################################
*/


`include "common.vh"

module sdram_init_loader #(parameter ROM_SIZE_IN_BYTES = (8 *1024))  (
    input wire                                      clk,
    input wire                                      reset_n,

    input  wire                                     dram_ack,
    output logic unsigned [`MEM_ADDR_BITS - 1 : 0]  dram_mem_addr,
    output logic                                    dram_mem_write_en,
    output wire  unsigned [`XLEN_BYTES - 1 : 0]     dram_mem_byte_enable,
    output logic unsigned [`XLEN - 1 : 0]           dram_mem_write_data,
    
    output logic                                    done
);

     logic [`XLEN - 1 : 0]                          rom_mem [0 : ROM_SIZE_IN_BYTES / 4 - 1];
     
     
     
     logic  unsigned [$clog2(ROM_SIZE_IN_BYTES / 4) - 1 : 0]    count;
     
     logic                                                      ctl_inc_count;
     logic                                                      ctl_load;
     
     
     always_ff @(posedge clk, negedge reset_n) begin
        if (!reset_n) begin
            count <= 0;
        end else if (ctl_inc_count) begin
            count <= count + 1;
        end
        
     end
     
     
     assign dram_mem_byte_enable = 4'b1111;
     
     always_ff @(posedge clk, negedge reset_n) begin
        if (!reset_n) begin
            dram_mem_write_en <= 0;
            dram_mem_addr <= 0;
            dram_mem_write_data <= 0;
        end else begin
            dram_mem_write_en <= ctl_load;
            dram_mem_addr <= count;
            dram_mem_write_data <= rom_mem[count];
        end
     end

    //+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
    // FSM
    //+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
        enum {S_IDLE, S_LOAD, S_WAIT, S_END} states;
                    
        localparam FSM_NUM_OF_STATES = states.num();
        logic [FSM_NUM_OF_STATES - 1:0] current_state = 0, next_state;
                    
        // Declare states
        always_ff @(posedge clk, negedge reset_n) begin : state_machine_reg
            if (!reset_n) begin
                current_state <= 0;
            end else begin
                current_state <= next_state;
            end
        end : state_machine_reg

        // state cast for debug, one-hot translation, enum value can be shown in the simulation in this way
        // Hopefully, synthesizer will optimize out the "states" variable

        // synthesis translate_off
        ///////////////////////////////////////////////////////////////////////
            always_comb begin : state_cast_for_debug
                for (int i = 0; i < FSM_NUM_OF_STATES; ++i) begin
                    if (current_state[i]) begin
                        $cast(states, i);
                    end
                end
            end : state_cast_for_debug
        ///////////////////////////////////////////////////////////////////////
        // synthesis translate_on   

        // FSM main body
        always_comb begin : state_machine_comb

            next_state = 0;
            
            ctl_inc_count = 0;
            ctl_load = 0;
            
            done = 0;
            
            case (1'b1) // synthesis parallel_case 

                current_state[S_IDLE]: begin
                    next_state [S_LOAD] = 1'b1;
                end

                current_state [S_LOAD] : begin
                    ctl_load = 1'b1;
                    next_state[S_WAIT] = 1'b1;

                end

                current_state [S_WAIT] : begin
                    if (dram_ack) begin
                        if (count == (ROM_SIZE_IN_BYTES /4 - 1)) begin
                            done = 1'b1;
                            next_state [S_END] = 1'b1;
                        end else begin
                            next_state[S_LOAD] = 1'b1;
                            ctl_inc_count = 1'b1;
                        end
                    end else begin
                        next_state [S_WAIT] = 1'b1;
                    end
                end
                
                current_state [S_END] : begin
                    next_state [S_END] = 1'b1;
                end
                
                default: begin
                    next_state[S_IDLE] = 1'b1;
                end

            endcase

        end : state_machine_comb  
     
     

//=================================================================================================================
// Initial data for ROM
//=================================================================================================================


initial begin

rom_mem[0] <= 32'h00003197;
rom_mem[1] <= 32'h55018193;
rom_mem[2] <= 32'h80818513;
rom_mem[3] <= 32'ha7c18613;
rom_mem[4] <= 32'h40a60633;
rom_mem[5] <= 32'h00000593;
rom_mem[6] <= 32'h3e0010ef;
rom_mem[7] <= 32'h00001517;
rom_mem[8] <= 32'h2e450513;
rom_mem[9] <= 32'h290010ef;
rom_mem[10] <= 32'h338010ef;
rom_mem[11] <= 32'h00012503;
rom_mem[12] <= 32'h00410593;
rom_mem[13] <= 32'h00000613;
rom_mem[14] <= 32'h0e0010ef;
rom_mem[15] <= 32'h28c0106f;
rom_mem[16] <= 32'h00008067;
rom_mem[17] <= 32'h00003517;
rom_mem[18] <= 32'hd0c50513;
rom_mem[19] <= 32'h00003797;
rom_mem[20] <= 32'hd0478793;
rom_mem[21] <= 32'h00a78a63;
rom_mem[22] <= 32'h80000317;
rom_mem[23] <= 32'hfa830313;
rom_mem[24] <= 32'h00030463;
rom_mem[25] <= 32'h00030067;
rom_mem[26] <= 32'h00008067;
rom_mem[27] <= 32'h00003517;
rom_mem[28] <= 32'hce450513;
rom_mem[29] <= 32'h00003597;
rom_mem[30] <= 32'hcdc58593;
rom_mem[31] <= 32'h40a585b3;
rom_mem[32] <= 32'h4025d593;
rom_mem[33] <= 32'h01f5d793;
rom_mem[34] <= 32'h00b785b3;
rom_mem[35] <= 32'h4015d593;
rom_mem[36] <= 32'h00058a63;
rom_mem[37] <= 32'h80000317;
rom_mem[38] <= 32'hf6c30313;
rom_mem[39] <= 32'h00030463;
rom_mem[40] <= 32'h00030067;
rom_mem[41] <= 32'h00008067;
rom_mem[42] <= 32'h8081c783;
rom_mem[43] <= 32'h04079063;
rom_mem[44] <= 32'hff010113;
rom_mem[45] <= 32'h00112623;
rom_mem[46] <= 32'hf8dff0ef;
rom_mem[47] <= 32'h80000797;
rom_mem[48] <= 32'hf4478793;
rom_mem[49] <= 32'h00078a63;
rom_mem[50] <= 32'h00002517;
rom_mem[51] <= 32'h83450513;
rom_mem[52] <= 32'h80000097;
rom_mem[53] <= 32'hf30080e7;
rom_mem[54] <= 32'h00c12083;
rom_mem[55] <= 32'h00100793;
rom_mem[56] <= 32'h80f18423;
rom_mem[57] <= 32'h01010113;
rom_mem[58] <= 32'h00008067;
rom_mem[59] <= 32'h00008067;
rom_mem[60] <= 32'h80000797;
rom_mem[61] <= 32'hf1078793;
rom_mem[62] <= 32'h02078663;
rom_mem[63] <= 32'hff010113;
rom_mem[64] <= 32'h83018593;
rom_mem[65] <= 32'h00001517;
rom_mem[66] <= 32'h7f850513;
rom_mem[67] <= 32'h00112623;
rom_mem[68] <= 32'h80000097;
rom_mem[69] <= 32'hef0080e7;
rom_mem[70] <= 32'h00c12083;
rom_mem[71] <= 32'h01010113;
rom_mem[72] <= 32'hf4dff06f;
rom_mem[73] <= 32'hf49ff06f;
rom_mem[74] <= 32'h200007b7;
rom_mem[75] <= 32'h0187c703;
rom_mem[76] <= 32'h01f77713;
rom_mem[77] <= 32'h02070063;
rom_mem[78] <= 32'h81118693;
rom_mem[79] <= 32'h0006c603;
rom_mem[80] <= 32'h00160793;
rom_mem[81] <= 32'h00f68023;
rom_mem[82] <= 32'h84818793;
rom_mem[83] <= 32'h00c787b3;
rom_mem[84] <= 32'h00e78023;
rom_mem[85] <= 32'h00008067;
rom_mem[86] <= 32'h300026f3;
rom_mem[87] <= 32'h30005073;
rom_mem[88] <= 32'h20000737;
rom_mem[89] <= 32'h00072783;
rom_mem[90] <= 32'h00472603;
rom_mem[91] <= 32'h00a78533;
rom_mem[92] <= 32'h00f537b3;
rom_mem[93] <= 32'h00c787b3;
rom_mem[94] <= 32'hfff00613;
rom_mem[95] <= 32'h00c72423;
rom_mem[96] <= 32'h00f72623;
rom_mem[97] <= 32'h00a72423;
rom_mem[98] <= 32'h30069073;
rom_mem[99] <= 32'h00008067;
rom_mem[100] <= 32'h81d1c703;
rom_mem[101] <= 32'h00100793;
rom_mem[102] <= 32'h200005b7;
rom_mem[103] <= 32'h00e797b3;
rom_mem[104] <= 32'h0ff7f793;
rom_mem[105] <= 32'h00f58ca3;
rom_mem[106] <= 32'h81d1c503;
rom_mem[107] <= 32'h81e1d703;
rom_mem[108] <= 32'h00251793;
rom_mem[109] <= 32'h80003637;
rom_mem[110] <= 32'h40f75733;
rom_mem[111] <= 32'h81c1c783;
rom_mem[112] <= 32'h00f77713;
rom_mem[113] <= 32'h91860613;
rom_mem[114] <= 32'h00c70733;
rom_mem[115] <= 32'h00074703;
rom_mem[116] <= 32'h40a7d7b3;
rom_mem[117] <= 32'h00779793;
rom_mem[118] <= 32'h00e7e7b3;
rom_mem[119] <= 32'h0ff7f793;
rom_mem[120] <= 32'h00f58c23;
rom_mem[121] <= 32'h81d1c783;
rom_mem[122] <= 32'h00178793;
rom_mem[123] <= 32'h0037f793;
rom_mem[124] <= 32'h80f18ea3;
rom_mem[125] <= 32'h8181a503;
rom_mem[126] <= 32'hf61ff06f;
rom_mem[127] <= 32'hfe010113;
rom_mem[128] <= 32'h00810693;
rom_mem[129] <= 32'h81418513;
rom_mem[130] <= 32'h00100713;
rom_mem[131] <= 32'h03000613;
rom_mem[132] <= 32'h05300593;
rom_mem[133] <= 32'h00112e23;
rom_mem[134] <= 32'h6c8000ef;
rom_mem[135] <= 32'h01c12083;
rom_mem[136] <= 32'h00814503;
rom_mem[137] <= 32'h02010113;
rom_mem[138] <= 32'h00008067;
rom_mem[139] <= 32'hfe010113;
rom_mem[140] <= 32'h00812c23;
rom_mem[141] <= 32'h00100713;
rom_mem[142] <= 32'h00f10693;
rom_mem[143] <= 32'h00000613;
rom_mem[144] <= 32'h05300593;
rom_mem[145] <= 32'h81418513;
rom_mem[146] <= 32'h00112e23;
rom_mem[147] <= 32'h694000ef;
rom_mem[148] <= 32'h00f14703;
rom_mem[149] <= 32'h0e500793;
rom_mem[150] <= 32'h00f70a63;
rom_mem[151] <= 32'h800015b7;
rom_mem[152] <= 32'h7b058593;
rom_mem[153] <= 32'ha4818513;
rom_mem[154] <= 32'h0f1000ef;
rom_mem[155] <= 32'h81418513;
rom_mem[156] <= 32'h00800693;
rom_mem[157] <= 32'h02d00613;
rom_mem[158] <= 32'h05300593;
rom_mem[159] <= 32'h5c4000ef;
rom_mem[160] <= 32'h81418513;
rom_mem[161] <= 32'h00600693;
rom_mem[162] <= 32'h02400613;
rom_mem[163] <= 32'h05300593;
rom_mem[164] <= 32'h5b0000ef;
rom_mem[165] <= 32'h81418513;
rom_mem[166] <= 32'h00300693;
rom_mem[167] <= 32'h02500613;
rom_mem[168] <= 32'h05300593;
rom_mem[169] <= 32'h59c000ef;
rom_mem[170] <= 32'h81418513;
rom_mem[171] <= 32'h00300693;
rom_mem[172] <= 32'h02600613;
rom_mem[173] <= 32'h05300593;
rom_mem[174] <= 32'h588000ef;
rom_mem[175] <= 32'h81418513;
rom_mem[176] <= 32'h0ff00693;
rom_mem[177] <= 32'h02700613;
rom_mem[178] <= 32'h05300593;
rom_mem[179] <= 32'h574000ef;
rom_mem[180] <= 32'h81418513;
rom_mem[181] <= 32'h00700693;
rom_mem[182] <= 32'h02c00613;
rom_mem[183] <= 32'h05300593;
rom_mem[184] <= 32'h560000ef;
rom_mem[185] <= 32'h81418513;
rom_mem[186] <= 32'h00000693;
rom_mem[187] <= 32'h02f00613;
rom_mem[188] <= 32'h05300593;
rom_mem[189] <= 32'h54c000ef;
rom_mem[190] <= 32'h81418513;
rom_mem[191] <= 32'h01000693;
rom_mem[192] <= 32'h02e00613;
rom_mem[193] <= 32'h05300593;
rom_mem[194] <= 32'h538000ef;
rom_mem[195] <= 32'h81418513;
rom_mem[196] <= 32'h00b00693;
rom_mem[197] <= 32'h03100613;
rom_mem[198] <= 32'h05300593;
rom_mem[199] <= 32'h524000ef;
rom_mem[200] <= 32'h81418513;
rom_mem[201] <= 32'h08000693;
rom_mem[202] <= 32'h03800613;
rom_mem[203] <= 32'h05300593;
rom_mem[204] <= 32'h510000ef;
rom_mem[205] <= 32'hec9ff0ef;
rom_mem[206] <= 32'h01c12083;
rom_mem[207] <= 32'h01812403;
rom_mem[208] <= 32'h02010113;
rom_mem[209] <= 32'h00008067;
rom_mem[210] <= 32'hfd010113;
rom_mem[211] <= 32'h03212023;
rom_mem[212] <= 32'h02812423;
rom_mem[213] <= 32'h02912223;
rom_mem[214] <= 32'h01312e23;
rom_mem[215] <= 32'h00100713;
rom_mem[216] <= 32'h00050993;
rom_mem[217] <= 32'h00058493;
rom_mem[218] <= 32'h00060413;
rom_mem[219] <= 32'h00710693;
rom_mem[220] <= 32'h00000613;
rom_mem[221] <= 32'h05300593;
rom_mem[222] <= 32'h81418513;
rom_mem[223] <= 32'h02112623;
rom_mem[224] <= 32'h560000ef;
rom_mem[225] <= 32'h00714703;
rom_mem[226] <= 32'h0e500793;
rom_mem[227] <= 32'h02f70463;
rom_mem[228] <= 32'h800015b7;
rom_mem[229] <= 32'h7b058593;
rom_mem[230] <= 32'ha4818513;
rom_mem[231] <= 32'h7bc000ef;
rom_mem[232] <= 32'h00714583;
rom_mem[233] <= 32'h01000613;
rom_mem[234] <= 32'ha4818513;
rom_mem[235] <= 32'h1b9000ef;
rom_mem[236] <= 32'h0000006f;
rom_mem[237] <= 32'he49ff0ef;
rom_mem[238] <= 32'h00a103a3;
rom_mem[239] <= 32'h01851513;
rom_mem[240] <= 32'h41855513;
rom_mem[241] <= 32'h08055a63;
rom_mem[242] <= 32'h00600713;
rom_mem[243] <= 32'h00810693;
rom_mem[244] <= 32'h03200613;
rom_mem[245] <= 32'h05300593;
rom_mem[246] <= 32'h81418513;
rom_mem[247] <= 32'h504000ef;
rom_mem[248] <= 32'h00914783;
rom_mem[249] <= 32'h00814703;
rom_mem[250] <= 32'h00879793;
rom_mem[251] <= 32'h00e7e7b3;
rom_mem[252] <= 32'h01379793;
rom_mem[253] <= 32'h0137d713;
rom_mem[254] <= 32'h0007d663;
rom_mem[255] <= 32'hffffe7b7;
rom_mem[256] <= 32'h00f76733;
rom_mem[257] <= 32'h00b14783;
rom_mem[258] <= 32'h00e99023;
rom_mem[259] <= 32'h00a14703;
rom_mem[260] <= 32'h00879793;
rom_mem[261] <= 32'h00e7e7b3;
rom_mem[262] <= 32'h01379793;
rom_mem[263] <= 32'h0137d713;
rom_mem[264] <= 32'h0007d663;
rom_mem[265] <= 32'hffffe7b7;
rom_mem[266] <= 32'h00f76733;
rom_mem[267] <= 32'h00d14783;
rom_mem[268] <= 32'h00e49023;
rom_mem[269] <= 32'h00c14703;
rom_mem[270] <= 32'h00879793;
rom_mem[271] <= 32'h00e7e7b3;
rom_mem[272] <= 32'h01379793;
rom_mem[273] <= 32'h0137d713;
rom_mem[274] <= 32'h0007d663;
rom_mem[275] <= 32'hffffe7b7;
rom_mem[276] <= 32'h00f76733;
rom_mem[277] <= 32'h00e41023;
rom_mem[278] <= 32'h00714783;
rom_mem[279] <= 32'h0107f793;
rom_mem[280] <= 32'h02078863;
rom_mem[281] <= 32'h800015b7;
rom_mem[282] <= 32'h7d458593;
rom_mem[283] <= 32'ha4818513;
rom_mem[284] <= 32'h6e8000ef;
rom_mem[285] <= 32'h800037b7;
rom_mem[286] <= 32'hd5078793;
rom_mem[287] <= 32'h0007c703;
rom_mem[288] <= 32'h200006b7;
rom_mem[289] <= 32'h00e68d23;
rom_mem[290] <= 32'hfff74713;
rom_mem[291] <= 32'h00e78023;
rom_mem[292] <= 32'h02c12083;
rom_mem[293] <= 32'h02812403;
rom_mem[294] <= 32'h00714503;
rom_mem[295] <= 32'h02412483;
rom_mem[296] <= 32'h02012903;
rom_mem[297] <= 32'h01c12983;
rom_mem[298] <= 32'h03010113;
rom_mem[299] <= 32'h00008067;
rom_mem[300] <= 32'hff010113;
rom_mem[301] <= 32'h3e800513;
rom_mem[302] <= 32'h00112623;
rom_mem[303] <= 32'h141000ef;
rom_mem[304] <= 32'hd6dff0ef;
rom_mem[305] <= 32'h8181a503;
rom_mem[306] <= 32'hc91ff0ef;
rom_mem[307] <= 32'h800005b7;
rom_mem[308] <= 32'h00300613;
rom_mem[309] <= 32'h19058593;
rom_mem[310] <= 32'h00000513;
rom_mem[311] <= 32'h33d000ef;
rom_mem[312] <= 32'h800015b7;
rom_mem[313] <= 32'h00300613;
rom_mem[314] <= 32'h80858593;
rom_mem[315] <= 32'h00100513;
rom_mem[316] <= 32'h329000ef;
rom_mem[317] <= 32'h800005b7;
rom_mem[318] <= 32'h00300613;
rom_mem[319] <= 32'h12858593;
rom_mem[320] <= 32'h01e00513;
rom_mem[321] <= 32'h315000ef;
rom_mem[322] <= 32'h0d5000ef;
rom_mem[323] <= 32'h1e300713;
rom_mem[324] <= 32'h00001537;
rom_mem[325] <= 32'h80e19f23;
rom_mem[326] <= 32'h38850513;
rom_mem[327] <= 32'h80018e23;
rom_mem[328] <= 32'h0dd000ef;
rom_mem[329] <= 32'h800037b7;
rom_mem[330] <= 32'h03f00713;
rom_mem[331] <= 32'h90e78c23;
rom_mem[332] <= 32'h91878793;
rom_mem[333] <= 32'h00600713;
rom_mem[334] <= 32'h00e780a3;
rom_mem[335] <= 32'h04f00713;
rom_mem[336] <= 32'h00e781a3;
rom_mem[337] <= 32'h00c12083;
rom_mem[338] <= 32'h01010113;
rom_mem[339] <= 32'h00008067;
rom_mem[340] <= 32'hfb010113;
rom_mem[341] <= 32'h05212023;
rom_mem[342] <= 32'h80c18793;
rom_mem[343] <= 32'h0007a583;
rom_mem[344] <= 32'h04812423;
rom_mem[345] <= 32'h04112623;
rom_mem[346] <= 32'h00a00613;
rom_mem[347] <= 32'h00158593;
rom_mem[348] <= 32'h04912223;
rom_mem[349] <= 32'h03312e23;
rom_mem[350] <= 32'h03412c23;
rom_mem[351] <= 32'h03512a23;
rom_mem[352] <= 32'h03612823;
rom_mem[353] <= 32'h03712623;
rom_mem[354] <= 32'h03812423;
rom_mem[355] <= 32'h03912223;
rom_mem[356] <= 32'h03a12023;
rom_mem[357] <= 32'h01b12e23;
rom_mem[358] <= 32'ha4818513;
rom_mem[359] <= 32'h00b7a023;
rom_mem[360] <= 32'h764000ef;
rom_mem[361] <= 32'h800015b7;
rom_mem[362] <= 32'h7e858593;
rom_mem[363] <= 32'ha4818513;
rom_mem[364] <= 32'h548000ef;
rom_mem[365] <= 32'h800015b7;
rom_mem[366] <= 32'h7ec58593;
rom_mem[367] <= 32'ha4818513;
rom_mem[368] <= 32'h538000ef;
rom_mem[369] <= 32'h200007b7;
rom_mem[370] <= 32'h0197c683;
rom_mem[371] <= 32'h00000593;
rom_mem[372] <= 32'h00000793;
rom_mem[373] <= 32'h0ff6f693;
rom_mem[374] <= 32'h80c18913;
rom_mem[375] <= 32'h00700813;
rom_mem[376] <= 32'h00800613;
rom_mem[377] <= 32'h40f6d733;
rom_mem[378] <= 32'h40f80533;
rom_mem[379] <= 32'h00177713;
rom_mem[380] <= 32'h00a71733;
rom_mem[381] <= 32'h00e585b3;
rom_mem[382] <= 32'h00178793;
rom_mem[383] <= 32'h0ff5f593;
rom_mem[384] <= 32'hfec792e3;
rom_mem[385] <= 32'h01000613;
rom_mem[386] <= 32'ha4818513;
rom_mem[387] <= 32'h754000ef;
rom_mem[388] <= 32'h800015b7;
rom_mem[389] <= 32'h7f458593;
rom_mem[390] <= 32'ha4818513;
rom_mem[391] <= 32'h4dc000ef;
rom_mem[392] <= 32'h8121c683;
rom_mem[393] <= 32'h8131c703;
rom_mem[394] <= 32'h81218493;
rom_mem[395] <= 32'h81318a13;
rom_mem[396] <= 32'h04e68863;
rom_mem[397] <= 32'h800025b7;
rom_mem[398] <= 32'h80458593;
rom_mem[399] <= 32'ha4818513;
rom_mem[400] <= 32'h4b8000ef;
rom_mem[401] <= 32'h94818993;
rom_mem[402] <= 32'h0004c583;
rom_mem[403] <= 32'h00100613;
rom_mem[404] <= 32'ha4818513;
rom_mem[405] <= 32'h00158793;
rom_mem[406] <= 32'h00b985b3;
rom_mem[407] <= 32'h00f48023;
rom_mem[408] <= 32'h3f4000ef;
rom_mem[409] <= 32'h0004c703;
rom_mem[410] <= 32'h000a4783;
rom_mem[411] <= 32'hfcf71ee3;
rom_mem[412] <= 32'h800025b7;
rom_mem[413] <= 32'h81458593;
rom_mem[414] <= 32'ha4818513;
rom_mem[415] <= 32'h47c000ef;
rom_mem[416] <= 32'h8101c703;
rom_mem[417] <= 32'h8111c783;
rom_mem[418] <= 32'h81018493;
rom_mem[419] <= 32'h81118993;
rom_mem[420] <= 32'h08f70c63;
rom_mem[421] <= 32'h800025b7;
rom_mem[422] <= 32'h81858593;
rom_mem[423] <= 32'ha4818513;
rom_mem[424] <= 32'h458000ef;
rom_mem[425] <= 32'h84818a13;
rom_mem[426] <= 32'h00100b13;
rom_mem[427] <= 32'h80002bb7;
rom_mem[428] <= 32'h80002c37;
rom_mem[429] <= 32'h80002cb7;
rom_mem[430] <= 32'h80002d37;
rom_mem[431] <= 32'h80002db7;
rom_mem[432] <= 32'h80002ab7;
rom_mem[433] <= 32'h0004c783;
rom_mem[434] <= 32'h828d8593;
rom_mem[435] <= 32'h00178713;
rom_mem[436] <= 32'h00fa07b3;
rom_mem[437] <= 32'h0007c783;
rom_mem[438] <= 32'h00e48023;
rom_mem[439] <= 32'h03678663;
rom_mem[440] <= 32'h00200713;
rom_mem[441] <= 32'h830d0593;
rom_mem[442] <= 32'h02e78063;
rom_mem[443] <= 32'h00400713;
rom_mem[444] <= 32'h838c8593;
rom_mem[445] <= 32'h00e78a63;
rom_mem[446] <= 32'h00800713;
rom_mem[447] <= 32'h840c0593;
rom_mem[448] <= 32'h00e78463;
rom_mem[449] <= 32'h844b8593;
rom_mem[450] <= 32'ha4818513;
rom_mem[451] <= 32'h44c000ef;
rom_mem[452] <= 32'h8aca8593;
rom_mem[453] <= 32'ha4818513;
rom_mem[454] <= 32'h440000ef;
rom_mem[455] <= 32'h0004c703;
rom_mem[456] <= 32'h0009c783;
rom_mem[457] <= 32'hfaf710e3;
rom_mem[458] <= 32'h00092703;
rom_mem[459] <= 32'h00e10613;
rom_mem[460] <= 32'h80e19f23;
rom_mem[461] <= 32'h00100713;
rom_mem[462] <= 32'h80e18e23;
rom_mem[463] <= 32'h20000737;
rom_mem[464] <= 32'hfff00793;
rom_mem[465] <= 32'h00f70d23;
rom_mem[466] <= 32'h01974783;
rom_mem[467] <= 32'h00c10593;
rom_mem[468] <= 32'h00a10513;
rom_mem[469] <= 32'hfff7c793;
rom_mem[470] <= 32'h0ff7f793;
rom_mem[471] <= 32'h00f70da3;
rom_mem[472] <= 32'hbe9ff0ef;
rom_mem[473] <= 32'h800025b7;
rom_mem[474] <= 32'h84c58593;
rom_mem[475] <= 32'ha4818513;
rom_mem[476] <= 32'h388000ef;
rom_mem[477] <= 32'h00a11583;
rom_mem[478] <= 32'h00a00613;
rom_mem[479] <= 32'ha4818513;
rom_mem[480] <= 32'h584000ef;
rom_mem[481] <= 32'h800025b7;
rom_mem[482] <= 32'h85458593;
rom_mem[483] <= 32'ha4818513;
rom_mem[484] <= 32'h368000ef;
rom_mem[485] <= 32'h00c11583;
rom_mem[486] <= 32'h00a00613;
rom_mem[487] <= 32'ha4818513;
rom_mem[488] <= 32'h564000ef;
rom_mem[489] <= 32'h800025b7;
rom_mem[490] <= 32'h85c58593;
rom_mem[491] <= 32'ha4818513;
rom_mem[492] <= 32'h348000ef;
rom_mem[493] <= 32'h00e11583;
rom_mem[494] <= 32'h00a00613;
rom_mem[495] <= 32'ha4818513;
rom_mem[496] <= 32'h548000ef;
rom_mem[497] <= 32'h3e800513;
rom_mem[498] <= 32'h634000ef;
rom_mem[499] <= 32'h04c12083;
rom_mem[500] <= 32'h04812403;
rom_mem[501] <= 32'h04412483;
rom_mem[502] <= 32'h04012903;
rom_mem[503] <= 32'h03c12983;
rom_mem[504] <= 32'h03812a03;
rom_mem[505] <= 32'h03412a83;
rom_mem[506] <= 32'h03012b03;
rom_mem[507] <= 32'h02c12b83;
rom_mem[508] <= 32'h02812c03;
rom_mem[509] <= 32'h02412c83;
rom_mem[510] <= 32'h02012d03;
rom_mem[511] <= 32'h01c12d83;
rom_mem[512] <= 32'h05010113;
rom_mem[513] <= 32'h00008067;
rom_mem[514] <= 32'hff010113;
rom_mem[515] <= 32'ha4818513;
rom_mem[516] <= 32'h00112623;
rom_mem[517] <= 32'h200000ef;
rom_mem[518] <= 32'h81318713;
rom_mem[519] <= 32'h00074683;
rom_mem[520] <= 32'h00168793;
rom_mem[521] <= 32'h00f70023;
rom_mem[522] <= 32'h94818793;
rom_mem[523] <= 32'h00d787b3;
rom_mem[524] <= 32'h00a78023;
rom_mem[525] <= 32'h00c12083;
rom_mem[526] <= 32'h01010113;
rom_mem[527] <= 32'h00008067;
rom_mem[528] <= 32'h200007b7;
rom_mem[529] <= 32'h00900713;
rom_mem[530] <= 32'h00159593;
rom_mem[531] <= 32'h02e78223;
rom_mem[532] <= 32'h0ff5f593;
rom_mem[533] <= 32'h0247c703;
rom_mem[534] <= 32'h02478513;
rom_mem[535] <= 32'h01871713;
rom_mem[536] <= 32'h41875713;
rom_mem[537] <= 32'hfe0758e3;
rom_mem[538] <= 32'h02b78423;
rom_mem[539] <= 32'h00a00793;
rom_mem[540] <= 32'h00f50023;
rom_mem[541] <= 32'h30005073;
rom_mem[542] <= 32'h20000737;
rom_mem[543] <= 32'h02474783;
rom_mem[544] <= 32'h0107f793;
rom_mem[545] <= 32'hfe078ce3;
rom_mem[546] <= 32'h02c70423;
rom_mem[547] <= 32'h20000737;
rom_mem[548] <= 32'h02474783;
rom_mem[549] <= 32'h0107f793;
rom_mem[550] <= 32'hfe078ce3;
rom_mem[551] <= 32'h02d70423;
rom_mem[552] <= 32'h200007b7;
rom_mem[553] <= 32'h0247c703;
rom_mem[554] <= 32'h02478693;
rom_mem[555] <= 32'h01077713;
rom_mem[556] <= 32'hfe070ae3;
rom_mem[557] <= 32'hfff00713;
rom_mem[558] <= 32'h02e78423;
rom_mem[559] <= 32'h30005073;
rom_mem[560] <= 32'h00800793;
rom_mem[561] <= 32'h00f68023;
rom_mem[562] <= 32'h20000737;
rom_mem[563] <= 32'h02474783;
rom_mem[564] <= 32'h01879793;
rom_mem[565] <= 32'h4187d793;
rom_mem[566] <= 32'hfe07dae3;
rom_mem[567] <= 32'h00008067;
rom_mem[568] <= 32'h30002873;
rom_mem[569] <= 32'h200007b7;
rom_mem[570] <= 32'h00900513;
rom_mem[571] <= 32'h00159593;
rom_mem[572] <= 32'h02a78223;
rom_mem[573] <= 32'h0ff5f593;
rom_mem[574] <= 32'h0247c503;
rom_mem[575] <= 32'h02478893;
rom_mem[576] <= 32'h01851513;
rom_mem[577] <= 32'h41855513;
rom_mem[578] <= 32'hfe0558e3;
rom_mem[579] <= 32'h02b78423;
rom_mem[580] <= 32'h00a00793;
rom_mem[581] <= 32'h00f88023;
rom_mem[582] <= 32'h30005073;
rom_mem[583] <= 32'h20000537;
rom_mem[584] <= 32'h02454783;
rom_mem[585] <= 32'h0107f793;
rom_mem[586] <= 32'hfe078ce3;
rom_mem[587] <= 32'h02c50423;
rom_mem[588] <= 32'h30081073;
rom_mem[589] <= 32'h200007b7;
rom_mem[590] <= 32'h0247c603;
rom_mem[591] <= 32'h02478513;
rom_mem[592] <= 32'h01067613;
rom_mem[593] <= 32'hfe060ae3;
rom_mem[594] <= 32'h02b78423;
rom_mem[595] <= 32'h01c00793;
rom_mem[596] <= 32'h00f50023;
rom_mem[597] <= 32'h20000637;
rom_mem[598] <= 32'h02464783;
rom_mem[599] <= 32'h01879793;
rom_mem[600] <= 32'h4187d793;
rom_mem[601] <= 32'hfe07dae3;
rom_mem[602] <= 32'h00e00793;
rom_mem[603] <= 32'h02f60223;
rom_mem[604] <= 32'h30005073;
rom_mem[605] <= 32'h00000793;
rom_mem[606] <= 32'h20000637;
rom_mem[607] <= 32'h0ff7f593;
rom_mem[608] <= 32'h02e5f463;
rom_mem[609] <= 32'h02464583;
rom_mem[610] <= 32'h0205f593;
rom_mem[611] <= 32'hfe058ce3;
rom_mem[612] <= 32'h02864503;
rom_mem[613] <= 32'h00f685b3;
rom_mem[614] <= 32'h00178793;
rom_mem[615] <= 32'h00a58023;
rom_mem[616] <= 32'h02060423;
rom_mem[617] <= 32'hfd9ff06f;
rom_mem[618] <= 32'h30081073;
rom_mem[619] <= 32'h00800713;
rom_mem[620] <= 32'h200007b7;
rom_mem[621] <= 32'h02e78223;
rom_mem[622] <= 32'h20000737;
rom_mem[623] <= 32'h02474783;
rom_mem[624] <= 32'h01879793;
rom_mem[625] <= 32'h4187d793;
rom_mem[626] <= 32'hfe07dae3;
rom_mem[627] <= 32'h00008067;
rom_mem[628] <= 32'hffffc7b7;
rom_mem[629] <= 32'heef78793;
rom_mem[630] <= 32'h80f19f23;
rom_mem[631] <= 32'h80018ea3;
rom_mem[632] <= 32'h80018e23;
rom_mem[633] <= 32'h000017b7;
rom_mem[634] <= 32'h9c478793;
rom_mem[635] <= 32'h80f1ac23;
rom_mem[636] <= 32'h00008067;
rom_mem[637] <= 32'h00008067;
rom_mem[638] <= 32'h200007b7;
rom_mem[639] <= 32'h0147a503;
rom_mem[640] <= 32'h01d55513;
rom_mem[641] <= 32'h00157513;
rom_mem[642] <= 32'h00008067;
rom_mem[643] <= 32'h00000513;
rom_mem[644] <= 32'h00008067;
rom_mem[645] <= 32'h200007b7;
rom_mem[646] <= 32'h80000737;
rom_mem[647] <= 32'h00e7aa23;
rom_mem[648] <= 32'h0147a503;
rom_mem[649] <= 32'h0ff57513;
rom_mem[650] <= 32'h00008067;
rom_mem[651] <= 32'h200007b7;
rom_mem[652] <= 32'h0107a683;
rom_mem[653] <= 32'hfe06cee3;
rom_mem[654] <= 32'h00b7a823;
rom_mem[655] <= 32'h00100513;
rom_mem[656] <= 32'h00008067;
rom_mem[657] <= 32'h200007b7;
rom_mem[658] <= 32'h10000737;
rom_mem[659] <= 32'h00e7aa23;
rom_mem[660] <= 32'h00008067;
rom_mem[661] <= 32'hfe010113;
rom_mem[662] <= 32'h00812c23;
rom_mem[663] <= 32'h00912a23;
rom_mem[664] <= 32'h01212823;
rom_mem[665] <= 32'h01312623;
rom_mem[666] <= 32'h00112e23;
rom_mem[667] <= 32'h00050913;
rom_mem[668] <= 32'h00058413;
rom_mem[669] <= 32'h00c589b3;
rom_mem[670] <= 32'h00000493;
rom_mem[671] <= 32'h03340263;
rom_mem[672] <= 32'h00092783;
rom_mem[673] <= 32'h00140413;
rom_mem[674] <= 32'hfff44583;
rom_mem[675] <= 32'h0007a783;
rom_mem[676] <= 32'h00090513;
rom_mem[677] <= 32'h000780e7;
rom_mem[678] <= 32'h00a484b3;
rom_mem[679] <= 32'hfe1ff06f;
rom_mem[680] <= 32'h01c12083;
rom_mem[681] <= 32'h01812403;
rom_mem[682] <= 32'h00048513;
rom_mem[683] <= 32'h01012903;
rom_mem[684] <= 32'h01412483;
rom_mem[685] <= 32'h00c12983;
rom_mem[686] <= 32'h02010113;
rom_mem[687] <= 32'h00008067;
rom_mem[688] <= 32'hfe010113;
rom_mem[689] <= 32'h00812c23;
rom_mem[690] <= 32'h00050413;
rom_mem[691] <= 32'h00058513;
rom_mem[692] <= 32'h00112e23;
rom_mem[693] <= 32'h00b12623;
rom_mem[694] <= 32'h1fd000ef;
rom_mem[695] <= 32'h00050613;
rom_mem[696] <= 32'h00040513;
rom_mem[697] <= 32'h01812403;
rom_mem[698] <= 32'h00c12583;
rom_mem[699] <= 32'h01c12083;
rom_mem[700] <= 32'h02010113;
rom_mem[701] <= 32'hf61ff06f;
rom_mem[702] <= 32'h00058463;
rom_mem[703] <= 32'hfc5ff06f;
rom_mem[704] <= 32'h00000513;
rom_mem[705] <= 32'h00008067;
rom_mem[706] <= 32'h00052783;
rom_mem[707] <= 32'h0007a303;
rom_mem[708] <= 32'h00030067;
rom_mem[709] <= 32'hff010113;
rom_mem[710] <= 32'h00d00593;
rom_mem[711] <= 32'h00112623;
rom_mem[712] <= 32'h00812423;
rom_mem[713] <= 32'h00912223;
rom_mem[714] <= 32'h00050493;
rom_mem[715] <= 32'hfddff0ef;
rom_mem[716] <= 32'h00050413;
rom_mem[717] <= 32'h00a00593;
rom_mem[718] <= 32'h00048513;
rom_mem[719] <= 32'hfcdff0ef;
rom_mem[720] <= 32'h00a40533;
rom_mem[721] <= 32'h00c12083;
rom_mem[722] <= 32'h00812403;
rom_mem[723] <= 32'h00412483;
rom_mem[724] <= 32'h01010113;
rom_mem[725] <= 32'h00008067;
rom_mem[726] <= 32'hff010113;
rom_mem[727] <= 32'h00812423;
rom_mem[728] <= 32'h00912223;
rom_mem[729] <= 32'h00112623;
rom_mem[730] <= 32'h00050493;
rom_mem[731] <= 32'h00000413;
rom_mem[732] <= 32'h00058663;
rom_mem[733] <= 32'hf4dff0ef;
rom_mem[734] <= 32'h00050413;
rom_mem[735] <= 32'h00048513;
rom_mem[736] <= 32'hf95ff0ef;
rom_mem[737] <= 32'h00850533;
rom_mem[738] <= 32'h00c12083;
rom_mem[739] <= 32'h00812403;
rom_mem[740] <= 32'h00412483;
rom_mem[741] <= 32'h01010113;
rom_mem[742] <= 32'h00008067;
rom_mem[743] <= 32'hfb010113;
rom_mem[744] <= 32'h04812423;
rom_mem[745] <= 32'h05212023;
rom_mem[746] <= 32'h03412c23;
rom_mem[747] <= 32'h04112623;
rom_mem[748] <= 32'h04912223;
rom_mem[749] <= 32'h03312e23;
rom_mem[750] <= 32'h03512a23;
rom_mem[751] <= 32'h02010623;
rom_mem[752] <= 32'h00100793;
rom_mem[753] <= 32'h00050a13;
rom_mem[754] <= 32'h00058913;
rom_mem[755] <= 32'h00a00413;
rom_mem[756] <= 32'h00c7f463;
rom_mem[757] <= 32'h00060413;
rom_mem[758] <= 32'h02c10493;
rom_mem[759] <= 32'h00900a93;
rom_mem[760] <= 32'h00040593;
rom_mem[761] <= 32'h00090513;
rom_mem[762] <= 32'h620000ef;
rom_mem[763] <= 32'h00050593;
rom_mem[764] <= 32'h00050993;
rom_mem[765] <= 32'h00040513;
rom_mem[766] <= 32'h554000ef;
rom_mem[767] <= 32'h40a90533;
rom_mem[768] <= 32'h0ff57513;
rom_mem[769] <= 32'h04aae863;
rom_mem[770] <= 32'h03050513;
rom_mem[771] <= 32'h0ff57513;
rom_mem[772] <= 32'hfff48493;
rom_mem[773] <= 32'h00a48023;
rom_mem[774] <= 32'h02897a63;
rom_mem[775] <= 32'h00048593;
rom_mem[776] <= 32'h000a0513;
rom_mem[777] <= 32'he9dff0ef;
rom_mem[778] <= 32'h04c12083;
rom_mem[779] <= 32'h04812403;
rom_mem[780] <= 32'h04412483;
rom_mem[781] <= 32'h04012903;
rom_mem[782] <= 32'h03c12983;
rom_mem[783] <= 32'h03812a03;
rom_mem[784] <= 32'h03412a83;
rom_mem[785] <= 32'h05010113;
rom_mem[786] <= 32'h00008067;
rom_mem[787] <= 32'h00098913;
rom_mem[788] <= 32'hf91ff06f;
rom_mem[789] <= 32'h03750513;
rom_mem[790] <= 32'hfb5ff06f;
rom_mem[791] <= 32'hff010113;
rom_mem[792] <= 32'h00812423;
rom_mem[793] <= 32'h00912223;
rom_mem[794] <= 32'h00112623;
rom_mem[795] <= 32'h01212023;
rom_mem[796] <= 32'h00050493;
rom_mem[797] <= 32'h00058413;
rom_mem[798] <= 32'h02061463;
rom_mem[799] <= 32'h00052703;
rom_mem[800] <= 32'h00812403;
rom_mem[801] <= 32'h00c12083;
rom_mem[802] <= 32'h00412483;
rom_mem[803] <= 32'h00012903;
rom_mem[804] <= 32'h00072303;
rom_mem[805] <= 32'h0ff5f593;
rom_mem[806] <= 32'h01010113;
rom_mem[807] <= 32'h00030067;
rom_mem[808] <= 32'h00a00813;
rom_mem[809] <= 32'h03061063;
rom_mem[810] <= 32'h0205c263;
rom_mem[811] <= 32'h00812403;
rom_mem[812] <= 32'h00c12083;
rom_mem[813] <= 32'h00412483;
rom_mem[814] <= 32'h00012903;
rom_mem[815] <= 32'h01010113;
rom_mem[816] <= 32'heddff06f;
rom_mem[817] <= 32'h0ff67613;
rom_mem[818] <= 32'hfe5ff06f;
rom_mem[819] <= 32'h02d00593;
rom_mem[820] <= 32'he39ff0ef;
rom_mem[821] <= 32'h00050913;
rom_mem[822] <= 32'h408005b3;
rom_mem[823] <= 32'h00048513;
rom_mem[824] <= 32'h00a00613;
rom_mem[825] <= 32'heb9ff0ef;
rom_mem[826] <= 32'h00c12083;
rom_mem[827] <= 32'h00812403;
rom_mem[828] <= 32'h00a90533;
rom_mem[829] <= 32'h00412483;
rom_mem[830] <= 32'h00012903;
rom_mem[831] <= 32'h01010113;
rom_mem[832] <= 32'h00008067;
rom_mem[833] <= 32'hf59ff06f;
rom_mem[834] <= 32'hff010113;
rom_mem[835] <= 32'h00112623;
rom_mem[836] <= 32'h00812423;
rom_mem[837] <= 32'h00912223;
rom_mem[838] <= 32'h00050493;
rom_mem[839] <= 32'hf41ff0ef;
rom_mem[840] <= 32'h00050413;
rom_mem[841] <= 32'h00048513;
rom_mem[842] <= 32'hdedff0ef;
rom_mem[843] <= 32'h00850533;
rom_mem[844] <= 32'h00c12083;
rom_mem[845] <= 32'h00812403;
rom_mem[846] <= 32'h00412483;
rom_mem[847] <= 32'h01010113;
rom_mem[848] <= 32'h00008067;
rom_mem[849] <= 32'h00061a63;
rom_mem[850] <= 32'h00052703;
rom_mem[851] <= 32'h0ff5f593;
rom_mem[852] <= 32'h00072303;
rom_mem[853] <= 32'h00030067;
rom_mem[854] <= 32'h0ff67613;
rom_mem[855] <= 32'he41ff06f;
rom_mem[856] <= 32'hfe5ff06f;
rom_mem[857] <= 32'hff010113;
rom_mem[858] <= 32'h00112623;
rom_mem[859] <= 32'h00812423;
rom_mem[860] <= 32'h00912223;
rom_mem[861] <= 32'h00050493;
rom_mem[862] <= 32'hfcdff0ef;
rom_mem[863] <= 32'h00050413;
rom_mem[864] <= 32'h00048513;
rom_mem[865] <= 32'hd91ff0ef;
rom_mem[866] <= 32'h00850533;
rom_mem[867] <= 32'h00c12083;
rom_mem[868] <= 32'h00812403;
rom_mem[869] <= 32'h00412483;
rom_mem[870] <= 32'h01010113;
rom_mem[871] <= 32'h00008067;
rom_mem[872] <= 32'hff010113;
rom_mem[873] <= 32'h00112623;
rom_mem[874] <= 32'h00812423;
rom_mem[875] <= 32'h00912223;
rom_mem[876] <= 32'h00050493;
rom_mem[877] <= 32'hf91ff0ef;
rom_mem[878] <= 32'h00050413;
rom_mem[879] <= 32'h00048513;
rom_mem[880] <= 32'hd55ff0ef;
rom_mem[881] <= 32'h00a40533;
rom_mem[882] <= 32'h00c12083;
rom_mem[883] <= 32'h00812403;
rom_mem[884] <= 32'h00412483;
rom_mem[885] <= 32'h01010113;
rom_mem[886] <= 32'h00008067;
rom_mem[887] <= 32'h000017b7;
rom_mem[888] <= 32'h88078793;
rom_mem[889] <= 32'h30479073;
rom_mem[890] <= 32'h30045073;
rom_mem[891] <= 32'h00008067;
rom_mem[892] <= 32'h30405073;
rom_mem[893] <= 32'h30005073;
rom_mem[894] <= 32'h00008067;
rom_mem[895] <= 32'hff010113;
rom_mem[896] <= 32'h00112623;
rom_mem[897] <= 32'h00812423;
rom_mem[898] <= 32'h00912223;
rom_mem[899] <= 32'h01212023;
rom_mem[900] <= 32'h30002973;
rom_mem[901] <= 32'h30005073;
rom_mem[902] <= 32'h200007b7;
rom_mem[903] <= 32'h0007a403;
rom_mem[904] <= 32'h0047a483;
rom_mem[905] <= 32'h30091073;
rom_mem[906] <= 32'h3e800613;
rom_mem[907] <= 32'h00000693;
rom_mem[908] <= 32'h00000593;
rom_mem[909] <= 32'h33c000ef;
rom_mem[910] <= 32'h00a40533;
rom_mem[911] <= 32'h00853433;
rom_mem[912] <= 32'h00b485b3;
rom_mem[913] <= 32'h00b405b3;
rom_mem[914] <= 32'h200007b7;
rom_mem[915] <= 32'h30005073;
rom_mem[916] <= 32'h0007a683;
rom_mem[917] <= 32'h0047a703;
rom_mem[918] <= 32'h30091073;
rom_mem[919] <= 32'hfeb768e3;
rom_mem[920] <= 32'h00e59463;
rom_mem[921] <= 32'hfea6e4e3;
rom_mem[922] <= 32'h00c12083;
rom_mem[923] <= 32'h00812403;
rom_mem[924] <= 32'h00412483;
rom_mem[925] <= 32'h00012903;
rom_mem[926] <= 32'h01010113;
rom_mem[927] <= 32'h00008067;
rom_mem[928] <= 32'ha4818793;
rom_mem[929] <= 32'h3e800713;
rom_mem[930] <= 32'h00e7a423;
rom_mem[931] <= 32'h80002737;
rom_mem[932] <= 32'h86c70713;
rom_mem[933] <= 32'h0007a223;
rom_mem[934] <= 32'h00e7a023;
rom_mem[935] <= 32'h00008067;
rom_mem[936] <= 32'hfb010113;
rom_mem[937] <= 32'h04112623;
rom_mem[938] <= 32'h04512423;
rom_mem[939] <= 32'h04612223;
rom_mem[940] <= 32'h04712023;
rom_mem[941] <= 32'h02812e23;
rom_mem[942] <= 32'h02912c23;
rom_mem[943] <= 32'h02a12a23;
rom_mem[944] <= 32'h02b12823;
rom_mem[945] <= 32'h02c12623;
rom_mem[946] <= 32'h02d12423;
rom_mem[947] <= 32'h02e12223;
rom_mem[948] <= 32'h02f12023;
rom_mem[949] <= 32'h01012e23;
rom_mem[950] <= 32'h01112c23;
rom_mem[951] <= 32'h01212a23;
rom_mem[952] <= 32'h01c12823;
rom_mem[953] <= 32'h01d12623;
rom_mem[954] <= 32'h01e12423;
rom_mem[955] <= 32'h01f12223;
rom_mem[956] <= 32'h342027f3;
rom_mem[957] <= 32'h0ff7f913;
rom_mem[958] <= 32'h300024f3;
rom_mem[959] <= 32'h30005073;
rom_mem[960] <= 32'h0807ce63;
rom_mem[961] <= 32'h800025b7;
rom_mem[962] <= 32'h8c858593;
rom_mem[963] <= 32'ha4818513;
rom_mem[964] <= 32'hbe9ff0ef;
rom_mem[965] <= 32'h01000613;
rom_mem[966] <= 32'h00090593;
rom_mem[967] <= 32'ha4818513;
rom_mem[968] <= 32'he45ff0ef;
rom_mem[969] <= 32'h800025b7;
rom_mem[970] <= 32'h8ec58593;
rom_mem[971] <= 32'ha4818513;
rom_mem[972] <= 32'hbc9ff0ef;
rom_mem[973] <= 32'h341025f3;
rom_mem[974] <= 32'h01000613;
rom_mem[975] <= 32'ha4818513;
rom_mem[976] <= 32'he61ff0ef;
rom_mem[977] <= 32'h30049073;
rom_mem[978] <= 32'h03c12403;
rom_mem[979] <= 32'h04c12083;
rom_mem[980] <= 32'h04812283;
rom_mem[981] <= 32'h04412303;
rom_mem[982] <= 32'h04012383;
rom_mem[983] <= 32'h03812483;
rom_mem[984] <= 32'h03412503;
rom_mem[985] <= 32'h03012583;
rom_mem[986] <= 32'h02c12603;
rom_mem[987] <= 32'h02812683;
rom_mem[988] <= 32'h02412703;
rom_mem[989] <= 32'h02012783;
rom_mem[990] <= 32'h01c12803;
rom_mem[991] <= 32'h01812883;
rom_mem[992] <= 32'h01412903;
rom_mem[993] <= 32'h01012e03;
rom_mem[994] <= 32'h00c12e83;
rom_mem[995] <= 32'h00812f03;
rom_mem[996] <= 32'h00412f83;
rom_mem[997] <= 32'h05010113;
rom_mem[998] <= 32'h30200073;
rom_mem[999] <= 32'h00700793;
rom_mem[1000] <= 32'h02f91063;
rom_mem[1001] <= 32'h344027f3;
rom_mem[1002] <= 32'hf7f7f793;
rom_mem[1003] <= 32'h34479073;
rom_mem[1004] <= 32'h82c1a783;
rom_mem[1005] <= 32'hf80788e3;
rom_mem[1006] <= 32'h000780e7;
rom_mem[1007] <= 32'hf89ff06f;
rom_mem[1008] <= 32'h200007b7;
rom_mem[1009] <= 32'h01c7a403;
rom_mem[1010] <= 32'h00247793;
rom_mem[1011] <= 32'h00078863;
rom_mem[1012] <= 32'h8201a783;
rom_mem[1013] <= 32'h00078463;
rom_mem[1014] <= 32'h000780e7;
rom_mem[1015] <= 32'h00141793;
rom_mem[1016] <= 32'h0007d863;
rom_mem[1017] <= 32'h8241a783;
rom_mem[1018] <= 32'h00078463;
rom_mem[1019] <= 32'h000780e7;
rom_mem[1020] <= 32'h00045863;
rom_mem[1021] <= 32'h8281a783;
rom_mem[1022] <= 32'h00078463;
rom_mem[1023] <= 32'h000780e7;
rom_mem[1024] <= 32'h344027f3;
rom_mem[1025] <= 32'hfffff737;
rom_mem[1026] <= 32'h7ff70713;
rom_mem[1027] <= 32'h00e7f7b3;
rom_mem[1028] <= 32'h34479073;
rom_mem[1029] <= 32'hf31ff06f;
rom_mem[1030] <= 32'hff010113;
rom_mem[1031] <= 32'h00112623;
rom_mem[1032] <= 32'h00812423;
rom_mem[1033] <= 32'h00912223;
rom_mem[1034] <= 32'h00300793;
rom_mem[1035] <= 32'h0af61463;
rom_mem[1036] <= 32'h00050413;
rom_mem[1037] <= 32'h00051e63;
rom_mem[1038] <= 32'h82b1a623;
rom_mem[1039] <= 32'h00c12083;
rom_mem[1040] <= 32'h00812403;
rom_mem[1041] <= 32'h00412483;
rom_mem[1042] <= 32'h01010113;
rom_mem[1043] <= 32'h00008067;
rom_mem[1044] <= 32'h00100513;
rom_mem[1045] <= 32'h00a41e63;
rom_mem[1046] <= 32'h20000737;
rom_mem[1047] <= 32'h82b1a023;
rom_mem[1048] <= 32'h02072783;
rom_mem[1049] <= 32'h0027e793;
rom_mem[1050] <= 32'h02f72023;
rom_mem[1051] <= 32'hfd1ff06f;
rom_mem[1052] <= 32'hfe240793;
rom_mem[1053] <= 32'h0ff7f713;
rom_mem[1054] <= 32'h02e56663;
rom_mem[1055] <= 32'h00279713;
rom_mem[1056] <= 32'h82418793;
rom_mem[1057] <= 32'h00e787b3;
rom_mem[1058] <= 32'h00b7a023;
rom_mem[1059] <= 32'h200007b7;
rom_mem[1060] <= 32'h0207a703;
rom_mem[1061] <= 32'h00851533;
rom_mem[1062] <= 32'h00e56533;
rom_mem[1063] <= 32'h02a7a023;
rom_mem[1064] <= 32'hf9dff06f;
rom_mem[1065] <= 32'h800025b7;
rom_mem[1066] <= 32'h88058593;
rom_mem[1067] <= 32'ha4818513;
rom_mem[1068] <= 32'ha49ff0ef;
rom_mem[1069] <= 32'h00040593;
rom_mem[1070] <= 32'h00812403;
rom_mem[1071] <= 32'h00c12083;
rom_mem[1072] <= 32'ha4818513;
rom_mem[1073] <= 32'h00412483;
rom_mem[1074] <= 32'h00a00613;
rom_mem[1075] <= 32'h01010113;
rom_mem[1076] <= 32'hc95ff06f;
rom_mem[1077] <= 32'h800025b7;
rom_mem[1078] <= 32'h89c58593;
rom_mem[1079] <= 32'ha4818513;
rom_mem[1080] <= 32'h00060493;
rom_mem[1081] <= 32'ha15ff0ef;
rom_mem[1082] <= 32'h00048593;
rom_mem[1083] <= 32'ha4818513;
rom_mem[1084] <= 32'h00a00613;
rom_mem[1085] <= 32'hc6dff0ef;
rom_mem[1086] <= 32'ha4818513;
rom_mem[1087] <= 32'h00812403;
rom_mem[1088] <= 32'h00c12083;
rom_mem[1089] <= 32'h00412483;
rom_mem[1090] <= 32'h800025b7;
rom_mem[1091] <= 32'h8b058593;
rom_mem[1092] <= 32'h01010113;
rom_mem[1093] <= 32'ha45ff06f;
rom_mem[1094] <= 32'hff010113;
rom_mem[1095] <= 32'h00112623;
rom_mem[1096] <= 32'hcd1ff0ef;
rom_mem[1097] <= 32'h0001c5b7;
rom_mem[1098] <= 32'h20058593;
rom_mem[1099] <= 32'ha4818513;
rom_mem[1100] <= 32'h915ff0ef;
rom_mem[1101] <= 32'h800017b7;
rom_mem[1102] <= 32'hea078793;
rom_mem[1103] <= 32'h30579073;
rom_mem[1104] <= 32'hb70ff0ef;
rom_mem[1105] <= 32'hc0cff0ef;
rom_mem[1106] <= 32'hffdff06f;
rom_mem[1107] <= 32'h00050613;
rom_mem[1108] <= 32'h00000513;
rom_mem[1109] <= 32'h0015f693;
rom_mem[1110] <= 32'h00068463;
rom_mem[1111] <= 32'h00c50533;
rom_mem[1112] <= 32'h0015d593;
rom_mem[1113] <= 32'h00161613;
rom_mem[1114] <= 32'hfe0596e3;
rom_mem[1115] <= 32'h00008067;
rom_mem[1116] <= 32'hff010113;
rom_mem[1117] <= 32'h00068293;
rom_mem[1118] <= 32'h00112623;
rom_mem[1119] <= 32'h00050393;
rom_mem[1120] <= 32'h00050693;
rom_mem[1121] <= 32'h00060713;
rom_mem[1122] <= 32'h00000793;
rom_mem[1123] <= 32'h00000313;
rom_mem[1124] <= 32'h00000813;
rom_mem[1125] <= 32'h010688b3;
rom_mem[1126] <= 32'h00177e93;
rom_mem[1127] <= 32'h00f30f33;
rom_mem[1128] <= 32'h01f6de13;
rom_mem[1129] <= 32'h00175713;
rom_mem[1130] <= 32'h0108bfb3;
rom_mem[1131] <= 32'h00179793;
rom_mem[1132] <= 32'h000e8663;
rom_mem[1133] <= 32'h01ef8333;
rom_mem[1134] <= 32'h00088813;
rom_mem[1135] <= 32'h00169693;
rom_mem[1136] <= 32'h01c7e7b3;
rom_mem[1137] <= 32'hfc0718e3;
rom_mem[1138] <= 32'h00058863;
rom_mem[1139] <= 32'h00060513;
rom_mem[1140] <= 32'hf7dff0ef;
rom_mem[1141] <= 32'h00a30333;
rom_mem[1142] <= 32'h00028a63;
rom_mem[1143] <= 32'h00038513;
rom_mem[1144] <= 32'h00028593;
rom_mem[1145] <= 32'hf69ff0ef;
rom_mem[1146] <= 32'h00650333;
rom_mem[1147] <= 32'h00c12083;
rom_mem[1148] <= 32'h00080513;
rom_mem[1149] <= 32'h00030593;
rom_mem[1150] <= 32'h01010113;
rom_mem[1151] <= 32'h00008067;
rom_mem[1152] <= 32'h06054063;
rom_mem[1153] <= 32'h0605c663;
rom_mem[1154] <= 32'h00058613;
rom_mem[1155] <= 32'h00050593;
rom_mem[1156] <= 32'hfff00513;
rom_mem[1157] <= 32'h02060c63;
rom_mem[1158] <= 32'h00100693;
rom_mem[1159] <= 32'h00b67a63;
rom_mem[1160] <= 32'h00c05863;
rom_mem[1161] <= 32'h00161613;
rom_mem[1162] <= 32'h00169693;
rom_mem[1163] <= 32'hfeb66ae3;
rom_mem[1164] <= 32'h00000513;
rom_mem[1165] <= 32'h00c5e663;
rom_mem[1166] <= 32'h40c585b3;
rom_mem[1167] <= 32'h00d56533;
rom_mem[1168] <= 32'h0016d693;
rom_mem[1169] <= 32'h00165613;
rom_mem[1170] <= 32'hfe0696e3;
rom_mem[1171] <= 32'h00008067;
rom_mem[1172] <= 32'h00008293;
rom_mem[1173] <= 32'hfb5ff0ef;
rom_mem[1174] <= 32'h00058513;
rom_mem[1175] <= 32'h00028067;
rom_mem[1176] <= 32'h40a00533;
rom_mem[1177] <= 32'h0005d863;
rom_mem[1178] <= 32'h40b005b3;
rom_mem[1179] <= 32'hf9dff06f;
rom_mem[1180] <= 32'h40b005b3;
rom_mem[1181] <= 32'h00008293;
rom_mem[1182] <= 32'hf91ff0ef;
rom_mem[1183] <= 32'h40a00533;
rom_mem[1184] <= 32'h00028067;
rom_mem[1185] <= 32'h00008293;
rom_mem[1186] <= 32'h0005ca63;
rom_mem[1187] <= 32'h00054c63;
rom_mem[1188] <= 32'hf79ff0ef;
rom_mem[1189] <= 32'h00058513;
rom_mem[1190] <= 32'h00028067;
rom_mem[1191] <= 32'h40b005b3;
rom_mem[1192] <= 32'hfe0558e3;
rom_mem[1193] <= 32'h40a00533;
rom_mem[1194] <= 32'hf61ff0ef;
rom_mem[1195] <= 32'h40b00533;
rom_mem[1196] <= 32'h00028067;
rom_mem[1197] <= 32'h00050593;
rom_mem[1198] <= 32'h00000693;
rom_mem[1199] <= 32'h00000613;
rom_mem[1200] <= 32'h00000513;
rom_mem[1201] <= 32'h29c0006f;
rom_mem[1202] <= 32'hff010113;
rom_mem[1203] <= 32'h00000593;
rom_mem[1204] <= 32'h00812423;
rom_mem[1205] <= 32'h00112623;
rom_mem[1206] <= 32'h00050413;
rom_mem[1207] <= 32'h390000ef;
rom_mem[1208] <= 32'h00000797;
rom_mem[1209] <= 32'h61878793;
rom_mem[1210] <= 32'h0007a503;
rom_mem[1211] <= 32'h03c52783;
rom_mem[1212] <= 32'h00078463;
rom_mem[1213] <= 32'h000780e7;
rom_mem[1214] <= 32'h00040513;
rom_mem[1215] <= 32'h4b0000ef;
rom_mem[1216] <= 32'hff010113;
rom_mem[1217] <= 32'h00812423;
rom_mem[1218] <= 32'h00001797;
rom_mem[1219] <= 32'h60878793;
rom_mem[1220] <= 32'h00001417;
rom_mem[1221] <= 32'h60440413;
rom_mem[1222] <= 32'h40f40433;
rom_mem[1223] <= 32'h00112623;
rom_mem[1224] <= 32'h00912223;
rom_mem[1225] <= 32'h40245413;
rom_mem[1226] <= 32'h02040263;
rom_mem[1227] <= 32'h00241493;
rom_mem[1228] <= 32'hffc48493;
rom_mem[1229] <= 32'h00f484b3;
rom_mem[1230] <= 32'h0004a783;
rom_mem[1231] <= 32'hfff40413;
rom_mem[1232] <= 32'hffc48493;
rom_mem[1233] <= 32'h000780e7;
rom_mem[1234] <= 32'hfe0418e3;
rom_mem[1235] <= 32'h00812403;
rom_mem[1236] <= 32'h00c12083;
rom_mem[1237] <= 32'h00412483;
rom_mem[1238] <= 32'h01010113;
rom_mem[1239] <= 32'hce5fe06f;
rom_mem[1240] <= 32'hff010113;
rom_mem[1241] <= 32'h00812423;
rom_mem[1242] <= 32'h01212023;
rom_mem[1243] <= 32'h00001417;
rom_mem[1244] <= 32'h59440413;
rom_mem[1245] <= 32'h00001917;
rom_mem[1246] <= 32'h58c90913;
rom_mem[1247] <= 32'h40890933;
rom_mem[1248] <= 32'h00112623;
rom_mem[1249] <= 32'h00912223;
rom_mem[1250] <= 32'h40295913;
rom_mem[1251] <= 32'h00090e63;
rom_mem[1252] <= 32'h00000493;
rom_mem[1253] <= 32'h00042783;
rom_mem[1254] <= 32'h00148493;
rom_mem[1255] <= 32'h00440413;
rom_mem[1256] <= 32'h000780e7;
rom_mem[1257] <= 32'hfe9918e3;
rom_mem[1258] <= 32'h00001417;
rom_mem[1259] <= 32'h55840413;
rom_mem[1260] <= 32'h00001917;
rom_mem[1261] <= 32'h56090913;
rom_mem[1262] <= 32'h40890933;
rom_mem[1263] <= 32'h40295913;
rom_mem[1264] <= 32'hc81fe0ef;
rom_mem[1265] <= 32'h00090e63;
rom_mem[1266] <= 32'h00000493;
rom_mem[1267] <= 32'h00042783;
rom_mem[1268] <= 32'h00148493;
rom_mem[1269] <= 32'h00440413;
rom_mem[1270] <= 32'h000780e7;
rom_mem[1271] <= 32'hfe9918e3;
rom_mem[1272] <= 32'h00c12083;
rom_mem[1273] <= 32'h00812403;
rom_mem[1274] <= 32'h00412483;
rom_mem[1275] <= 32'h00012903;
rom_mem[1276] <= 32'h01010113;
rom_mem[1277] <= 32'h00008067;
rom_mem[1278] <= 32'h00f00313;
rom_mem[1279] <= 32'h00050713;
rom_mem[1280] <= 32'h02c37e63;
rom_mem[1281] <= 32'h00f77793;
rom_mem[1282] <= 32'h0a079063;
rom_mem[1283] <= 32'h08059263;
rom_mem[1284] <= 32'hff067693;
rom_mem[1285] <= 32'h00f67613;
rom_mem[1286] <= 32'h00e686b3;
rom_mem[1287] <= 32'h00b72023;
rom_mem[1288] <= 32'h00b72223;
rom_mem[1289] <= 32'h00b72423;
rom_mem[1290] <= 32'h00b72623;
rom_mem[1291] <= 32'h01070713;
rom_mem[1292] <= 32'hfed766e3;
rom_mem[1293] <= 32'h00061463;
rom_mem[1294] <= 32'h00008067;
rom_mem[1295] <= 32'h40c306b3;
rom_mem[1296] <= 32'h00269693;
rom_mem[1297] <= 32'h00000297;
rom_mem[1298] <= 32'h005686b3;
rom_mem[1299] <= 32'h00c68067;
rom_mem[1300] <= 32'h00b70723;
rom_mem[1301] <= 32'h00b706a3;
rom_mem[1302] <= 32'h00b70623;
rom_mem[1303] <= 32'h00b705a3;
rom_mem[1304] <= 32'h00b70523;
rom_mem[1305] <= 32'h00b704a3;
rom_mem[1306] <= 32'h00b70423;
rom_mem[1307] <= 32'h00b703a3;
rom_mem[1308] <= 32'h00b70323;
rom_mem[1309] <= 32'h00b702a3;
rom_mem[1310] <= 32'h00b70223;
rom_mem[1311] <= 32'h00b701a3;
rom_mem[1312] <= 32'h00b70123;
rom_mem[1313] <= 32'h00b700a3;
rom_mem[1314] <= 32'h00b70023;
rom_mem[1315] <= 32'h00008067;
rom_mem[1316] <= 32'h0ff5f593;
rom_mem[1317] <= 32'h00859693;
rom_mem[1318] <= 32'h00d5e5b3;
rom_mem[1319] <= 32'h01059693;
rom_mem[1320] <= 32'h00d5e5b3;
rom_mem[1321] <= 32'hf6dff06f;
rom_mem[1322] <= 32'h00279693;
rom_mem[1323] <= 32'h00000297;
rom_mem[1324] <= 32'h005686b3;
rom_mem[1325] <= 32'h00008293;
rom_mem[1326] <= 32'hfa0680e7;
rom_mem[1327] <= 32'h00028093;
rom_mem[1328] <= 32'hff078793;
rom_mem[1329] <= 32'h40f70733;
rom_mem[1330] <= 32'h00f60633;
rom_mem[1331] <= 32'hf6c378e3;
rom_mem[1332] <= 32'hf3dff06f;
rom_mem[1333] <= 32'h00357793;
rom_mem[1334] <= 32'h00050713;
rom_mem[1335] <= 32'h04079c63;
rom_mem[1336] <= 32'h7f7f86b7;
rom_mem[1337] <= 32'hf7f68693;
rom_mem[1338] <= 32'hfff00593;
rom_mem[1339] <= 32'h00470713;
rom_mem[1340] <= 32'hffc72603;
rom_mem[1341] <= 32'h00d677b3;
rom_mem[1342] <= 32'h00d787b3;
rom_mem[1343] <= 32'h00c7e7b3;
rom_mem[1344] <= 32'h00d7e7b3;
rom_mem[1345] <= 32'hfeb784e3;
rom_mem[1346] <= 32'hffc74683;
rom_mem[1347] <= 32'h40a707b3;
rom_mem[1348] <= 32'hffd74603;
rom_mem[1349] <= 32'hffe74503;
rom_mem[1350] <= 32'h04068063;
rom_mem[1351] <= 32'h02060a63;
rom_mem[1352] <= 32'h00a03533;
rom_mem[1353] <= 32'h00f50533;
rom_mem[1354] <= 32'hffe50513;
rom_mem[1355] <= 32'h00008067;
rom_mem[1356] <= 32'hfa0688e3;
rom_mem[1357] <= 32'h00074783;
rom_mem[1358] <= 32'h00170713;
rom_mem[1359] <= 32'h00377693;
rom_mem[1360] <= 32'hfe0798e3;
rom_mem[1361] <= 32'h40a70733;
rom_mem[1362] <= 32'hfff70513;
rom_mem[1363] <= 32'h00008067;
rom_mem[1364] <= 32'hffd78513;
rom_mem[1365] <= 32'h00008067;
rom_mem[1366] <= 32'hffc78513;
rom_mem[1367] <= 32'h00008067;
rom_mem[1368] <= 32'hfe010113;
rom_mem[1369] <= 32'h00812c23;
rom_mem[1370] <= 32'h00001417;
rom_mem[1371] <= 32'h7ec40413;
rom_mem[1372] <= 32'h00912a23;
rom_mem[1373] <= 32'h00050493;
rom_mem[1374] <= 32'h00042503;
rom_mem[1375] <= 32'h01212823;
rom_mem[1376] <= 32'h01312623;
rom_mem[1377] <= 32'h01412423;
rom_mem[1378] <= 32'h00112e23;
rom_mem[1379] <= 32'h00058913;
rom_mem[1380] <= 32'h00060a13;
rom_mem[1381] <= 32'h00068993;
rom_mem[1382] <= 32'h20c000ef;
rom_mem[1383] <= 32'h00000797;
rom_mem[1384] <= 32'h35c78793;
rom_mem[1385] <= 32'h0007a703;
rom_mem[1386] <= 32'h14872783;
rom_mem[1387] <= 32'h08078663;
rom_mem[1388] <= 32'h0047a703;
rom_mem[1389] <= 32'h01f00813;
rom_mem[1390] <= 32'h00042503;
rom_mem[1391] <= 32'h08e84463;
rom_mem[1392] <= 32'h00271813;
rom_mem[1393] <= 32'h02049e63;
rom_mem[1394] <= 32'h00170713;
rom_mem[1395] <= 32'h00e7a223;
rom_mem[1396] <= 32'h010787b3;
rom_mem[1397] <= 32'h0127a423;
rom_mem[1398] <= 32'h1d0000ef;
rom_mem[1399] <= 32'h00000513;
rom_mem[1400] <= 32'h01c12083;
rom_mem[1401] <= 32'h01812403;
rom_mem[1402] <= 32'h01412483;
rom_mem[1403] <= 32'h01012903;
rom_mem[1404] <= 32'h00c12983;
rom_mem[1405] <= 32'h00812a03;
rom_mem[1406] <= 32'h02010113;
rom_mem[1407] <= 32'h00008067;
rom_mem[1408] <= 32'h010785b3;
rom_mem[1409] <= 32'h0945a423;
rom_mem[1410] <= 32'h1887a683;
rom_mem[1411] <= 32'h00100613;
rom_mem[1412] <= 32'h00e61633;
rom_mem[1413] <= 32'h00c6e6b3;
rom_mem[1414] <= 32'h18d7a423;
rom_mem[1415] <= 32'h1135a423;
rom_mem[1416] <= 32'h00200693;
rom_mem[1417] <= 32'hfad492e3;
rom_mem[1418] <= 32'h18c7a683;
rom_mem[1419] <= 32'h00c6e633;
rom_mem[1420] <= 32'h18c7a623;
rom_mem[1421] <= 32'hf95ff06f;
rom_mem[1422] <= 32'h14c70793;
rom_mem[1423] <= 32'h14f72423;
rom_mem[1424] <= 32'hf71ff06f;
rom_mem[1425] <= 32'h164000ef;
rom_mem[1426] <= 32'hfff00513;
rom_mem[1427] <= 32'hf95ff06f;
rom_mem[1428] <= 32'h7ffff797;
rom_mem[1429] <= 32'h9b078793;
rom_mem[1430] <= 32'h00078863;
rom_mem[1431] <= 32'h00000517;
rom_mem[1432] <= 32'hca450513;
rom_mem[1433] <= 32'hc51ff06f;
rom_mem[1434] <= 32'h00008067;
rom_mem[1435] <= 32'hfd010113;
rom_mem[1436] <= 32'h01612823;
rom_mem[1437] <= 32'h80418b13;
rom_mem[1438] <= 32'h01512a23;
rom_mem[1439] <= 32'h00050a93;
rom_mem[1440] <= 32'h000b2503;
rom_mem[1441] <= 32'h01312e23;
rom_mem[1442] <= 32'h01412c23;
rom_mem[1443] <= 32'h01712623;
rom_mem[1444] <= 32'h01912223;
rom_mem[1445] <= 32'h02112623;
rom_mem[1446] <= 32'h02812423;
rom_mem[1447] <= 32'h02912223;
rom_mem[1448] <= 32'h03212023;
rom_mem[1449] <= 32'h01812423;
rom_mem[1450] <= 32'h00058b93;
rom_mem[1451] <= 32'h0f8000ef;
rom_mem[1452] <= 32'h00000797;
rom_mem[1453] <= 32'h24878793;
rom_mem[1454] <= 32'h0007ac83;
rom_mem[1455] <= 32'h00100a13;
rom_mem[1456] <= 32'hfff00993;
rom_mem[1457] <= 32'h148ca903;
rom_mem[1458] <= 32'h02090863;
rom_mem[1459] <= 32'h00492483;
rom_mem[1460] <= 32'hfff48413;
rom_mem[1461] <= 32'h02044263;
rom_mem[1462] <= 32'h00249493;
rom_mem[1463] <= 32'h009904b3;
rom_mem[1464] <= 32'h040b8863;
rom_mem[1465] <= 32'h1044a783;
rom_mem[1466] <= 32'h05778463;
rom_mem[1467] <= 32'hfff40413;
rom_mem[1468] <= 32'hffc48493;
rom_mem[1469] <= 32'hff3416e3;
rom_mem[1470] <= 32'h02812403;
rom_mem[1471] <= 32'h000b2503;
rom_mem[1472] <= 32'h02c12083;
rom_mem[1473] <= 32'h02412483;
rom_mem[1474] <= 32'h02012903;
rom_mem[1475] <= 32'h01c12983;
rom_mem[1476] <= 32'h01812a03;
rom_mem[1477] <= 32'h01412a83;
rom_mem[1478] <= 32'h01012b03;
rom_mem[1479] <= 32'h00c12b83;
rom_mem[1480] <= 32'h00812c03;
rom_mem[1481] <= 32'h00412c83;
rom_mem[1482] <= 32'h03010113;
rom_mem[1483] <= 32'h07c0006f;
rom_mem[1484] <= 32'h00492783;
rom_mem[1485] <= 32'h0044a683;
rom_mem[1486] <= 32'hfff78793;
rom_mem[1487] <= 32'h04878a63;
rom_mem[1488] <= 32'h0004a223;
rom_mem[1489] <= 32'hfa0684e3;
rom_mem[1490] <= 32'h18892783;
rom_mem[1491] <= 32'h008a1733;
rom_mem[1492] <= 32'h00492c03;
rom_mem[1493] <= 32'h00f777b3;
rom_mem[1494] <= 32'h00079e63;
rom_mem[1495] <= 32'h000680e7;
rom_mem[1496] <= 32'h00492783;
rom_mem[1497] <= 32'hf78790e3;
rom_mem[1498] <= 32'h148ca783;
rom_mem[1499] <= 32'hf92780e3;
rom_mem[1500] <= 32'hf55ff06f;
rom_mem[1501] <= 32'h18c92783;
rom_mem[1502] <= 32'h0844a583;
rom_mem[1503] <= 32'h00f77733;
rom_mem[1504] <= 32'h00071c63;
rom_mem[1505] <= 32'h000a8513;
rom_mem[1506] <= 32'h000680e7;
rom_mem[1507] <= 32'hfd5ff06f;
rom_mem[1508] <= 32'h00892223;
rom_mem[1509] <= 32'hfb1ff06f;
rom_mem[1510] <= 32'h00058513;
rom_mem[1511] <= 32'h000680e7;
rom_mem[1512] <= 32'hfc1ff06f;
rom_mem[1513] <= 32'h00008067;
rom_mem[1514] <= 32'h00008067;
rom_mem[1515] <= 32'h0000006f;
rom_mem[1516] <= 32'h4c584441;
rom_mem[1517] <= 32'h20353433;
rom_mem[1518] <= 32'h69766564;
rom_mem[1519] <= 32'h49206563;
rom_mem[1520] <= 32'h6e752044;
rom_mem[1521] <= 32'h6f636572;
rom_mem[1522] <= 32'h7a696e67;
rom_mem[1523] <= 32'h21216465;
rom_mem[1524] <= 32'h00212121;
rom_mem[1525] <= 32'h4c445841;
rom_mem[1526] <= 32'h20353433;
rom_mem[1527] <= 32'h49544341;
rom_mem[1528] <= 32'h59544956;
rom_mem[1529] <= 32'h00000000;
rom_mem[1530] <= 32'h0000203a;
rom_mem[1531] <= 32'h3d205753;
rom_mem[1532] <= 32'h00783020;
rom_mem[1533] <= 32'h3d3d3d20;
rom_mem[1534] <= 32'h3d3d3d3d;
rom_mem[1535] <= 32'h203d3d3d;
rom_mem[1536] <= 32'h00000000;
rom_mem[1537] <= 32'h6f47200a;
rom_mem[1538] <= 32'h654d2074;
rom_mem[1539] <= 32'h67617373;
rom_mem[1540] <= 32'h00203a65;
rom_mem[1541] <= 32'h0000000a;
rom_mem[1542] <= 32'h654b200a;
rom_mem[1543] <= 32'h72502079;
rom_mem[1544] <= 32'h65737365;
rom_mem[1545] <= 32'h00203a64;
rom_mem[1546] <= 32'h66654c20;
rom_mem[1547] <= 32'h00000074;
rom_mem[1548] <= 32'h6e654320;
rom_mem[1549] <= 32'h00726574;
rom_mem[1550] <= 32'h776f4420;
rom_mem[1551] <= 32'h0000006e;
rom_mem[1552] <= 32'h00705520;
rom_mem[1553] <= 32'h67695220;
rom_mem[1554] <= 32'h00007468;
rom_mem[1555] <= 32'h203d2058;
rom_mem[1556] <= 32'h00000000;
rom_mem[1557] <= 32'h2059202c;
rom_mem[1558] <= 32'h0000203d;
rom_mem[1559] <= 32'h205a202c;
rom_mem[1560] <= 32'h0000203d;
rom_mem[1561] <= 32'h00000000;
rom_mem[1562] <= 32'h00000000;
rom_mem[1563] <= 32'h80000a2c;
rom_mem[1564] <= 32'h800009f8;
rom_mem[1565] <= 32'h80000a14;
rom_mem[1566] <= 32'h80000a0c;
rom_mem[1567] <= 32'h800009f4;
rom_mem[1568] <= 32'h6e6b6e75;
rom_mem[1569] <= 32'h206e776f;
rom_mem[1570] <= 32'h65746e69;
rom_mem[1571] <= 32'h70757272;
rom_mem[1572] <= 32'h6e692074;
rom_mem[1573] <= 32'h20786564;
rom_mem[1574] <= 32'h00000000;
rom_mem[1575] <= 32'h75736e75;
rom_mem[1576] <= 32'h726f7070;
rom_mem[1577] <= 32'h20646574;
rom_mem[1578] <= 32'h65646f6d;
rom_mem[1579] <= 32'h00000020;
rom_mem[1580] <= 32'h726f6620;
rom_mem[1581] <= 32'h74746120;
rom_mem[1582] <= 32'h49686361;
rom_mem[1583] <= 32'h7265746e;
rom_mem[1584] <= 32'h74707572;
rom_mem[1585] <= 32'h00000000;
rom_mem[1586] <= 32'h65637845;
rom_mem[1587] <= 32'h6f697470;
rom_mem[1588] <= 32'h2121206e;
rom_mem[1589] <= 32'h20212121;
rom_mem[1590] <= 32'h65637845;
rom_mem[1591] <= 32'h6f697470;
rom_mem[1592] <= 32'h6f43206e;
rom_mem[1593] <= 32'h3d206564;
rom_mem[1594] <= 32'h00783020;
rom_mem[1595] <= 32'h4350454d;
rom_mem[1596] <= 32'h30203d20;
rom_mem[1597] <= 32'h00000078;
rom_mem[1598] <= 32'h80002928;
rom_mem[1599] <= 32'h00000000;
rom_mem[2624] <= 32'h80001650;
rom_mem[2625] <= 32'h800000f0;
rom_mem[2626] <= 32'h800009d0;
rom_mem[2627] <= 32'h80000e80;
rom_mem[2628] <= 32'h800000a8;
rom_mem[2630] <= 32'h735b786d;
rom_mem[2631] <= 32'h077d6d66;
rom_mem[2632] <= 32'h7c776f7f;
rom_mem[2633] <= 32'h71795e39;
rom_mem[2634] <= 32'h00000000;
rom_mem[2635] <= 32'h80002c14;
rom_mem[2636] <= 32'h80002c7c;
rom_mem[2637] <= 32'h80002ce4;
rom_mem[2638] <= 32'h00000000;
rom_mem[2639] <= 32'h00000000;
rom_mem[2640] <= 32'h00000000;
rom_mem[2641] <= 32'h00000000;
rom_mem[2642] <= 32'h00000000;
rom_mem[2643] <= 32'h00000000;
rom_mem[2644] <= 32'h00000000;
rom_mem[2645] <= 32'h00000000;
rom_mem[2646] <= 32'h00000000;
rom_mem[2647] <= 32'h00000000;
rom_mem[2648] <= 32'h00000000;
rom_mem[2649] <= 32'h00000000;
rom_mem[2650] <= 32'h00000000;
rom_mem[2651] <= 32'h00000000;
rom_mem[2652] <= 32'h00000000;
rom_mem[2653] <= 32'h00000000;
rom_mem[2654] <= 32'h00000000;
rom_mem[2655] <= 32'h00000000;
rom_mem[2656] <= 32'h00000000;
rom_mem[2657] <= 32'h00000000;
rom_mem[2658] <= 32'h00000000;
rom_mem[2659] <= 32'h00000000;
rom_mem[2660] <= 32'h00000000;
rom_mem[2661] <= 32'h00000000;
rom_mem[2662] <= 32'h00000000;
rom_mem[2663] <= 32'h00000000;
rom_mem[2664] <= 32'h00000000;
rom_mem[2665] <= 32'h00000000;
rom_mem[2666] <= 32'h00000000;
rom_mem[2667] <= 32'h00000000;
rom_mem[2668] <= 32'h00000000;
rom_mem[2669] <= 32'h00000000;
rom_mem[2670] <= 32'h00000000;
rom_mem[2671] <= 32'h00000000;
rom_mem[2672] <= 32'h00000000;
rom_mem[2673] <= 32'h00000000;
rom_mem[2674] <= 32'h00000000;
rom_mem[2675] <= 32'h00000000;
rom_mem[2676] <= 32'h00000001;
rom_mem[2677] <= 32'h00000000;
rom_mem[2678] <= 32'habcd330e;
rom_mem[2679] <= 32'he66d1234;
rom_mem[2680] <= 32'h0005deec;
rom_mem[2681] <= 32'h0000000b;
rom_mem[2682] <= 32'h00000000;
rom_mem[2683] <= 32'h00000000;
rom_mem[2684] <= 32'h00000000;
rom_mem[2685] <= 32'h00000000;
rom_mem[2686] <= 32'h00000000;
rom_mem[2687] <= 32'h00000000;
rom_mem[2688] <= 32'h00000000;
rom_mem[2689] <= 32'h00000000;
rom_mem[2690] <= 32'h00000000;
rom_mem[2691] <= 32'h00000000;
rom_mem[2692] <= 32'h00000000;
rom_mem[2693] <= 32'h00000000;
rom_mem[2694] <= 32'h00000000;
rom_mem[2695] <= 32'h00000000;
rom_mem[2696] <= 32'h00000000;
rom_mem[2697] <= 32'h00000000;
rom_mem[2698] <= 32'h00000000;
rom_mem[2699] <= 32'h00000000;
rom_mem[2700] <= 32'h00000000;
rom_mem[2701] <= 32'h00000000;
rom_mem[2702] <= 32'h00000000;
rom_mem[2703] <= 32'h00000000;
rom_mem[2704] <= 32'h00000000;
rom_mem[2705] <= 32'h00000000;
rom_mem[2706] <= 32'h00000000;
rom_mem[2707] <= 32'h00000000;
rom_mem[2708] <= 32'h00000000;
rom_mem[2709] <= 32'h00000000;
rom_mem[2710] <= 32'h00000000;
rom_mem[2711] <= 32'h00000000;
rom_mem[2712] <= 32'h00000000;
rom_mem[2713] <= 32'h00000000;
rom_mem[2714] <= 32'h00000000;
rom_mem[2715] <= 32'h00000000;
rom_mem[2716] <= 32'h00000000;
rom_mem[2717] <= 32'h00000000;
rom_mem[2718] <= 32'h00000000;
rom_mem[2719] <= 32'h00000000;
rom_mem[2720] <= 32'h00000000;
rom_mem[2721] <= 32'h00000000;
rom_mem[2722] <= 32'h00000000;
rom_mem[2723] <= 32'h00000000;
rom_mem[2724] <= 32'h00000000;
rom_mem[2725] <= 32'h00000000;
rom_mem[2726] <= 32'h00000000;
rom_mem[2727] <= 32'h00000000;
rom_mem[2728] <= 32'h00000000;
rom_mem[2729] <= 32'h00000000;
rom_mem[2730] <= 32'h00000000;
rom_mem[2731] <= 32'h00000000;
rom_mem[2732] <= 32'h00000000;
rom_mem[2733] <= 32'h00000000;
rom_mem[2734] <= 32'h00000000;
rom_mem[2735] <= 32'h00000000;
rom_mem[2736] <= 32'h00000000;
rom_mem[2737] <= 32'h00000000;
rom_mem[2738] <= 32'h00000000;
rom_mem[2739] <= 32'h00000000;
rom_mem[2740] <= 32'h00000000;
rom_mem[2741] <= 32'h00000000;
rom_mem[2742] <= 32'h00000000;
rom_mem[2743] <= 32'h00000000;
rom_mem[2744] <= 32'h00000000;
rom_mem[2745] <= 32'h00000000;
rom_mem[2746] <= 32'h00000000;
rom_mem[2747] <= 32'h00000000;
rom_mem[2748] <= 32'h00000000;
rom_mem[2749] <= 32'h00000000;
rom_mem[2750] <= 32'h00000000;
rom_mem[2751] <= 32'h00000000;
rom_mem[2752] <= 32'h00000000;
rom_mem[2753] <= 32'h00000000;
rom_mem[2754] <= 32'h00000000;
rom_mem[2755] <= 32'h00000000;
rom_mem[2756] <= 32'h00000000;
rom_mem[2757] <= 32'h00000000;
rom_mem[2758] <= 32'h00000000;
rom_mem[2759] <= 32'h00000000;
rom_mem[2760] <= 32'h00000000;
rom_mem[2761] <= 32'h00000000;
rom_mem[2762] <= 32'h00000000;
rom_mem[2763] <= 32'h00000000;
rom_mem[2764] <= 32'h00000000;
rom_mem[2765] <= 32'h00000000;
rom_mem[2766] <= 32'h00000000;
rom_mem[2767] <= 32'h00000000;
rom_mem[2768] <= 32'h00000000;
rom_mem[2769] <= 32'h00000000;
rom_mem[2770] <= 32'h00000000;
rom_mem[2771] <= 32'h00000000;
rom_mem[2772] <= 32'h00000000;
rom_mem[2773] <= 32'h00000000;
rom_mem[2774] <= 32'h00000000;
rom_mem[2775] <= 32'h00000000;
rom_mem[2776] <= 32'h00000000;
rom_mem[2777] <= 32'h00000000;
rom_mem[2778] <= 32'h00000000;
rom_mem[2779] <= 32'h00000000;
rom_mem[2780] <= 32'h00000000;
rom_mem[2781] <= 32'h00000000;
rom_mem[2782] <= 32'h00000000;
rom_mem[2783] <= 32'h00000000;
rom_mem[2784] <= 32'h00000000;
rom_mem[2785] <= 32'h00000000;
rom_mem[2786] <= 32'h00000000;
rom_mem[2787] <= 32'h00000000;
rom_mem[2788] <= 32'h00000000;
rom_mem[2789] <= 32'h00000000;
rom_mem[2790] <= 32'h00000000;
rom_mem[2791] <= 32'h00000000;
rom_mem[2792] <= 32'h00000000;
rom_mem[2793] <= 32'h00000000;
rom_mem[2794] <= 32'h00000000;
rom_mem[2795] <= 32'h00000000;
rom_mem[2796] <= 32'h00000000;
rom_mem[2797] <= 32'h00000000;
rom_mem[2798] <= 32'h00000000;
rom_mem[2799] <= 32'h00000000;
rom_mem[2800] <= 32'h00000000;
rom_mem[2801] <= 32'h00000000;
rom_mem[2802] <= 32'h00000000;
rom_mem[2803] <= 32'h00000000;
rom_mem[2804] <= 32'h00000000;
rom_mem[2805] <= 32'h00000000;
rom_mem[2806] <= 32'h00000000;
rom_mem[2807] <= 32'h00000000;
rom_mem[2808] <= 32'h00000000;
rom_mem[2809] <= 32'h00000000;
rom_mem[2810] <= 32'h00000000;
rom_mem[2811] <= 32'h00000000;
rom_mem[2812] <= 32'h00000000;
rom_mem[2813] <= 32'h00000000;
rom_mem[2814] <= 32'h00000000;
rom_mem[2815] <= 32'h00000000;
rom_mem[2816] <= 32'h00000000;
rom_mem[2817] <= 32'h00000000;
rom_mem[2818] <= 32'h00000000;
rom_mem[2819] <= 32'h00000000;
rom_mem[2820] <= 32'h00000000;
rom_mem[2821] <= 32'h00000000;
rom_mem[2822] <= 32'h00000000;
rom_mem[2823] <= 32'h00000000;
rom_mem[2824] <= 32'h00000000;
rom_mem[2825] <= 32'h00000000;
rom_mem[2826] <= 32'h00000000;
rom_mem[2827] <= 32'h00000000;
rom_mem[2828] <= 32'h00000000;
rom_mem[2829] <= 32'h00000000;
rom_mem[2830] <= 32'h00000000;
rom_mem[2831] <= 32'h00000000;
rom_mem[2832] <= 32'h00000000;
rom_mem[2833] <= 32'h00000000;
rom_mem[2834] <= 32'h00000000;
rom_mem[2835] <= 32'h00000000;
rom_mem[2836] <= 32'h00000000;
rom_mem[2837] <= 32'h00000000;
rom_mem[2838] <= 32'h00000000;
rom_mem[2839] <= 32'h00000000;
rom_mem[2840] <= 32'h00000000;
rom_mem[2841] <= 32'h00000000;
rom_mem[2842] <= 32'h00000000;
rom_mem[2843] <= 32'h00000000;
rom_mem[2844] <= 32'h00000000;
rom_mem[2845] <= 32'h00000000;
rom_mem[2846] <= 32'h00000000;
rom_mem[2847] <= 32'h00000000;
rom_mem[2848] <= 32'h00000000;
rom_mem[2849] <= 32'h00000000;
rom_mem[2850] <= 32'h00000000;
rom_mem[2851] <= 32'h00000000;
rom_mem[2852] <= 32'h00000000;
rom_mem[2853] <= 32'h00000000;
rom_mem[2854] <= 32'h00000000;
rom_mem[2855] <= 32'h00000000;
rom_mem[2856] <= 32'h00000000;
rom_mem[2857] <= 32'h00000000;
rom_mem[2858] <= 32'h00000000;
rom_mem[2859] <= 32'h00000000;
rom_mem[2860] <= 32'h00000000;
rom_mem[2861] <= 32'h00000000;
rom_mem[2862] <= 32'h00000000;
rom_mem[2863] <= 32'h00000000;
rom_mem[2864] <= 32'h00000000;
rom_mem[2865] <= 32'h00000000;
rom_mem[2866] <= 32'h00000000;
rom_mem[2867] <= 32'h00000000;
rom_mem[2868] <= 32'h00000000;
rom_mem[2869] <= 32'h00000000;
rom_mem[2870] <= 32'h00000000;
rom_mem[2871] <= 32'h00000000;
rom_mem[2872] <= 32'h00000000;
rom_mem[2873] <= 32'h00000000;
rom_mem[2874] <= 32'h00000000;
rom_mem[2875] <= 32'h00000000;
rom_mem[2876] <= 32'h00000000;
rom_mem[2877] <= 32'h00000000;
rom_mem[2878] <= 32'h00000000;
rom_mem[2879] <= 32'h00000000;
rom_mem[2880] <= 32'h00000000;
rom_mem[2881] <= 32'h00000000;
rom_mem[2882] <= 32'h00000000;
rom_mem[2883] <= 32'h00000000;
rom_mem[2884] <= 32'h00000000;
rom_mem[2885] <= 32'h00000000;
rom_mem[2886] <= 32'h00000000;
rom_mem[2887] <= 32'h00000000;
rom_mem[2888] <= 32'h00000000;
rom_mem[2889] <= 32'h00000000;
rom_mem[2890] <= 32'h00000000;
rom_mem[2891] <= 32'h00000000;
rom_mem[2892] <= 32'h00000000;
rom_mem[2893] <= 32'h00000000;
rom_mem[2894] <= 32'h00000000;
rom_mem[2895] <= 32'h00000000;
rom_mem[2896] <= 32'h00000000;
rom_mem[2897] <= 32'h00000000;
rom_mem[2898] <= 32'h00000000;
rom_mem[2899] <= 32'h00000000;
rom_mem[2900] <= 32'h0000005a;
rom_mem[2901] <= 32'h80002fa8;

end

endmodule



