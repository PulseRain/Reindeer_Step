// ocd.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module ocd (
		input  wire         acq_clk,        // acq_clk.clk
		input  wire [255:0] acq_data_in,    //     tap.acq_data_in
		input  wire [3:0]   acq_trigger_in  //        .acq_trigger_in
	);

	sld_signaltap #(
		.sld_data_bits               (256),
		.sld_sample_depth            (1024),
		.sld_ram_block_type          ("AUTO"),
		.sld_storage_qualifier_mode  ("OFF"),
		.sld_trigger_bits            (4),
		.sld_trigger_level           (1),
		.sld_trigger_in_enabled      (0),
		.sld_enable_advanced_trigger (0),
		.sld_trigger_level_pipeline  (1),
		.sld_trigger_pipeline        (0),
		.sld_ram_pipeline            (0),
		.sld_counter_pipeline        (0),
		.sld_node_info               (806383104),
		.sld_incremental_routing     (0),
		.sld_node_crc_bits           (32),
		.sld_node_crc_hiword         (8522),
		.sld_node_crc_loword         (55810)
	) signaltap_ii_logic_analyzer_0 (
		.acq_data_in    (acq_data_in),    //     tap.acq_data_in
		.acq_trigger_in (acq_trigger_in), //        .acq_trigger_in
		.acq_clk        (acq_clk)         // acq_clk.clk
	);

endmodule
